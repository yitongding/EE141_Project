`include "Opcode.vh"
`include "const.vh"

module controller(
    input wire  [:0] datapath_contents,
    output wire [:0]  dpath_controls_i,
    output wire [:0]  exec_controls_x,
    output wire [:0]   hazard_controls
);


endmodule
