/**
 * UC Berkeley CS150
 * Fall 2014
 * List of ALU operations.
<<<<<<< HEAD
 */

=======
*/
>>>>>>> ca6419d66242e2742bb6de10b8f8c6853efdd5e3
`ifndef ALUOP
`define ALUOP

`define ALU_ADD     4'd0
`define ALU_SUB     4'd1
`define ALU_AND     4'd2
`define ALU_OR      4'd3
`define ALU_XOR     4'd4
`define ALU_SLT     4'd5
`define ALU_SLTU    4'd6
`define ALU_SLL     4'd7
`define ALU_SRA     4'd8
`define ALU_SRL     4'd9
`define ALU_COPY_B  4'd10
`define ALU_JALR    4'd11
`define ALU_XXX     4'd15

`endif //ALUOP
